
module f_box (
  input  logic [7:0] iword,
  output logic [7:0] oword
);


always @(*) begin
    case(iword)
      8'h00: oword = 8'hA3;
      8'h01: oword = 8'hD7;
      8'h02: oword = 8'h09;
      8'h03: oword = 8'h83;
      8'h04: oword = 8'hF8;
      8'h05: oword = 8'h48;
      8'h06: oword = 8'hF6;
      8'h07: oword = 8'hF4;
      8'h08: oword = 8'hB3;
      8'h09: oword = 8'h21;
      8'h0A: oword = 8'h15;
      8'h0B: oword = 8'h78;
      8'h0C: oword = 8'h99;
      8'h0D: oword = 8'hB1;
      8'h0E: oword = 8'hAF;
      8'h0F: oword = 8'hF9;
      8'h10: oword = 8'hE7;
      8'h11: oword = 8'h2D;
      8'h12: oword = 8'h4D;
      8'h13: oword = 8'h8A;
      8'h14: oword = 8'hCE;
      8'h15: oword = 8'h4C;
      8'h16: oword = 8'hCA;
      8'h17: oword = 8'h2E;
      8'h18: oword = 8'h52;
      8'h19: oword = 8'h95;
      8'h1A: oword = 8'hD9;
      8'h1B: oword = 8'h1E;
      8'h1C: oword = 8'h4E;
      8'h1D: oword = 8'h38;
      8'h1E: oword = 8'h44;
      8'h1F: oword = 8'h28;
      8'h20: oword = 8'h0A;
      8'h21: oword = 8'hDF;
      8'h22: oword = 8'h02;
      8'h23: oword = 8'hA0;
      8'h24: oword = 8'h17;
      8'h25: oword = 8'hF1;
      8'h26: oword = 8'h60;
      8'h27: oword = 8'h68;
      8'h28: oword = 8'h12;
      8'h29: oword = 8'hB7;
      8'h2A: oword = 8'h7A;
      8'h2B: oword = 8'hC3;
      8'h2C: oword = 8'hC9;
      8'h2D: oword = 8'hFA;
      8'h2E: oword = 8'h3D;
      8'h2F: oword = 8'h53;
      8'h30: oword = 8'h96;
      8'h31: oword = 8'h84;
      8'h32: oword = 8'h6B;
      8'h33: oword = 8'hBA;
      8'h34: oword = 8'hF2;
      8'h35: oword = 8'h63;
      8'h36: oword = 8'h9A;
      8'h37: oword = 8'h19;
      8'h38: oword = 8'h7C;
      8'h39: oword = 8'hAE;
      8'h3A: oword = 8'hE5;
      8'h3B: oword = 8'hF5;
      8'h3C: oword = 8'hF7;
      8'h3D: oword = 8'h16;
      8'h3E: oword = 8'h6A;
      8'h3F: oword = 8'hA2;
      8'h40: oword = 8'h39;
      8'h41: oword = 8'hB6;
      8'h42: oword = 8'h7B;
      8'h43: oword = 8'h0F;
      8'h44: oword = 8'hC1;
      8'h45: oword = 8'h93;
      8'h46: oword = 8'h81;
      8'h47: oword = 8'h1B;
      8'h48: oword = 8'hEE;
      8'h49: oword = 8'hB4;
      8'h4A: oword = 8'h1A;
      8'h4B: oword = 8'hEA;
      8'h4C: oword = 8'hD0;
      8'h4D: oword = 8'h91;
      8'h4E: oword = 8'h2F;
      8'h4F: oword = 8'hB8;
      8'h50: oword = 8'h55;
      8'h51: oword = 8'hB9;
      8'h52: oword = 8'hDA;
      8'h53: oword = 8'h85;
      8'h54: oword = 8'h3F;
      8'h55: oword = 8'h41;
      8'h56: oword = 8'hBF;
      8'h57: oword = 8'hE0;
      8'h58: oword = 8'h5A;
      8'h59: oword = 8'h58;
      8'h5A: oword = 8'h80;
      8'h5B: oword = 8'h5F;
      8'h5C: oword = 8'h66;
      8'h5D: oword = 8'h0B;
      8'h5E: oword = 8'hD8;
      8'h5F: oword = 8'h90;
      8'h60: oword = 8'h35;
      8'h61: oword = 8'hD5;
      8'h62: oword = 8'hC0;
      8'h63: oword = 8'hA7;
      8'h64: oword = 8'h33;
      8'h65: oword = 8'h06;
      8'h66: oword = 8'h65;
      8'h67: oword = 8'h69;
      8'h68: oword = 8'h45;
      8'h69: oword = 8'h00;
      8'h6A: oword = 8'h94;
      8'h6B: oword = 8'h56;
      8'h6C: oword = 8'h6D;
      8'h6D: oword = 8'h98;
      8'h6E: oword = 8'h9B;
      8'h6F: oword = 8'h76;
      8'h70: oword = 8'h97;
      8'h71: oword = 8'hFC;
      8'h72: oword = 8'hB2;
      8'h73: oword = 8'hC2;
      8'h74: oword = 8'hB0;
      8'h75: oword = 8'hFE;
      8'h76: oword = 8'hDB;
      8'h77: oword = 8'h20;
      8'h78: oword = 8'hE1;
      8'h79: oword = 8'hEB;
      8'h7A: oword = 8'hD6;
      8'h7B: oword = 8'hE4;
      8'h7C: oword = 8'hDD;
      8'h7D: oword = 8'h47;
      8'h7E: oword = 8'h4A;
      8'h7F: oword = 8'h1D;
      8'h80: oword = 8'h42;
      8'h81: oword = 8'hED;
      8'h82: oword = 8'h9E;
      8'h83: oword = 8'h6E;
      8'h84: oword = 8'h49;
      8'h85: oword = 8'h3C;
      8'h86: oword = 8'hCD;
      8'h87: oword = 8'h43;
      8'h88: oword = 8'h27;
      8'h89: oword = 8'hD2;
      8'h8A: oword = 8'h07;
      8'h8B: oword = 8'hD4;
      8'h8C: oword = 8'hDE;
      8'h8D: oword = 8'hC7;
      8'h8E: oword = 8'h67;
      8'h8F: oword = 8'h18;
      8'h90: oword = 8'h89;
      8'h91: oword = 8'hCB;
      8'h92: oword = 8'h30;
      8'h93: oword = 8'h1F;
      8'h94: oword = 8'h8D;
      8'h95: oword = 8'hC6;
      8'h96: oword = 8'h8F;
      8'h97: oword = 8'hAA;
      8'h98: oword = 8'hC8;
      8'h99: oword = 8'h74;
      8'h9A: oword = 8'hDC;
      8'h9B: oword = 8'hC9;
      8'h9C: oword = 8'h5D;
      8'h9D: oword = 8'h5C;
      8'h9E: oword = 8'h31;
      8'h9F: oword = 8'hA4;
      8'hA0: oword = 8'h70;
      8'hA1: oword = 8'h88;
      8'hA2: oword = 8'h61;
      8'hA3: oword = 8'h2C;
      8'hA4: oword = 8'h9F;
      8'hA5: oword = 8'h0D;
      8'hA6: oword = 8'h2B;
      8'hA7: oword = 8'h87;
      8'hA8: oword = 8'h50;
      8'hA9: oword = 8'h82;
      8'hAA: oword = 8'h54;
      8'hAB: oword = 8'h64;
      8'hAC: oword = 8'h26;
      8'hAD: oword = 8'h7D;
      8'hAE: oword = 8'h03;
      8'hAF: oword = 8'h40;
      8'hB0: oword = 8'h34;
      8'hB1: oword = 8'h4B;
      8'hB2: oword = 8'h1C;
      8'hB3: oword = 8'h73;
      8'hB4: oword = 8'hD1;
      8'hB5: oword = 8'hC4;
      8'hB6: oword = 8'hFD;
      8'hB7: oword = 8'h3B;
      8'hB8: oword = 8'hCC;
      8'hB9: oword = 8'hFB;
      8'hBA: oword = 8'h7F;
      8'hBB: oword = 8'hAB;
      8'hBC: oword = 8'hE6;
      8'hBD: oword = 8'h3E;
      8'hBE: oword = 8'h5B;
      8'hBF: oword = 8'hA5;
      8'hC0: oword = 8'hAD;
      8'hC1: oword = 8'h04;
      8'hC2: oword = 8'h23;
      8'hC3: oword = 8'h9C;
      8'hC4: oword = 8'h14;
      8'hC5: oword = 8'h51;
      8'hC6: oword = 8'h22;
      8'hC7: oword = 8'hF0;
      8'hC8: oword = 8'h29;
      8'hC9: oword = 8'h79;
      8'hCA: oword = 8'h71;
      8'hCB: oword = 8'h7E;
      8'hCC: oword = 8'hFF;
      8'hCD: oword = 8'h8C;
      8'hCE: oword = 8'h0E;
      8'hCF: oword = 8'hE2;
      8'hD0: oword = 8'h0C;
      8'hD1: oword = 8'hEF;
      8'hD2: oword = 8'hBC;
      8'hD3: oword = 8'h72;
      8'hD4: oword = 8'h75;
      8'hD5: oword = 8'h6F;
      8'hD6: oword = 8'h37;
      8'hD7: oword = 8'hA1;
      8'hD8: oword = 8'hEC;
      8'hD9: oword = 8'hD3;
      8'hDA: oword = 8'h8E;
      8'hDB: oword = 8'h62;
      8'hDC: oword = 8'h8B;
      8'hDD: oword = 8'h86;
      8'hDE: oword = 8'h10;
      8'hDF: oword = 8'hE8;
      8'hE0: oword = 8'h08;
      8'hE1: oword = 8'h77;
      8'hE2: oword = 8'h11;
      8'hE3: oword = 8'hBE;
      8'hE4: oword = 8'h92;
      8'hE5: oword = 8'h4F;
      8'hE6: oword = 8'h24;
      8'hE7: oword = 8'hC5;
      8'hE8: oword = 8'h32;
      8'hE9: oword = 8'h36;
      8'hEA: oword = 8'h9D;
      8'hEB: oword = 8'hCF;
      8'hEC: oword = 8'hF3;
      8'hED: oword = 8'hA6;
      8'hEE: oword = 8'hBB;
      8'hEF: oword = 8'hAC;
      8'hF0: oword = 8'h5E;
      8'hF1: oword = 8'h6C;
      8'hF2: oword = 8'hA9;
      8'hF3: oword = 8'h13;
      8'hF4: oword = 8'h57;
      8'hF5: oword = 8'h25;
      8'hF6: oword = 8'hB5;
      8'hF7: oword = 8'hE3;
      8'hF8: oword = 8'hBD;
      8'hF9: oword = 8'hA8;
      8'hFA: oword = 8'h3A;
      8'hFB: oword = 8'h01;
      8'hFC: oword = 8'h05;
      8'hFD: oword = 8'h59;
      8'hFE: oword = 8'h2A;
      8'hFF: oword = 8'h46;
    endcase
  end

endmodule